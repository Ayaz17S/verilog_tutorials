module or_gate(f,x,y);
input x,y;
output f;
assign f = x|y;
endmodule